library ieee;
use ieee.std_logic_1164.all;

entity control_fast is
	port (	-- Input
			clk : in std_logic;
			reset : in std_logic;
			opcode : in std_logic_vector(5 downto 0);
			-- Output 
			pc_write_cond : out std_logic;
			pc_write : out std_logic;
			i_or_d : out std_logic;
			mem_read : out std_logic;
			mem_write : out std_logic;
			mem_to_reg : out std_logic;
			ir_write : out std_logic;
			reg_dest : out std_logic;
			reg_write : out std_logic;
			alu_src_a : out std_logic;
			alu_src_b : out std_logic_vector(1 downto 0);
			alu_op : out std_logic_vector(1 downto 0);
			pc_source : out std_logic_vector(1 downto 0));	
end entity;

architecture fsm of control_fast is		 

type state_type is (
	inst_fetch, 
	inst_decode_reg_fetch,
	execution,
	r_comp,
	mem_comp,  
	branch_comp, 
	jump_comp, 
	mem_w, 
	mem_r, 
	write_back);

attribute enum_encoding : string;
attribute enum_encoding of
state_type : type is "0000 0001 0011 0010 1000 1001 0101 1010 1100 0100";
	
signal current_state : state_type; 

begin			  
	
	control_output : process (current_state, opcode)
	begin
		
		pc_write_cond <= '0';
		pc_write <= '0'; 
		i_or_d <= '0'; 
		mem_read <= '0'; 
		mem_write <= '0';
		mem_to_reg <= '0'; 
		ir_write <= '0';
		reg_dest <= '0'; 
		reg_write <= '0'; 
		alu_src_a <= '0'; 
		alu_src_b <= "00";
		alu_op <= "00";
		pc_source <= "00";
		
		case current_state is
			when inst_fetch => 
				pc_write <= '1'; 
				i_or_d <= '0'; 
				mem_read <= '1'; 
				ir_write <= '1';
				-- alu_src_a <= '0'; 
				alu_src_b <= "00";
				alu_op <= "00";
				pc_source <= "00";
			when inst_decode_reg_fetch =>  
				-- alu_src_a <= '0'; 
				alu_src_b <= "00";
				-- alu_op <= '00';
			when mem_comp =>	 
				alu_src_a <= '1'; 
				alu_src_b <= "00";
				-- alu_op <= '00';
			when execution => 
				alu_src_a <= '1'; 
				-- alu_src_b <= '00';
				alu_op <= "00";
			when branch_comp => 
				pc_write_cond <= '1';
				alu_src_a <= '1'; 
				-- alu_src_b <= '00';
				alu_op <= "00";
				pc_source <= "00";
			when jump_comp => 
				pc_write <= '1'; 
				pc_source <= "00";
			when mem_r => 
				i_or_d <= '1'; 
				mem_read <= '1'; 	
			when mem_w => 
				i_or_d <= '1'; 
				mem_write <= '1';
			when r_comp =>
				-- mem_to_reg <= '0'; 
				reg_dest <= '1'; 
				reg_write <= '1'; 
			when write_back => 
				mem_to_reg <= '1'; 
				reg_dest <= '1'; 
				reg_write <= '1';
			when others =>
				null;
		end case;
	end process;
	
	fsm_state : process (clk, reset)
	begin		
		if reset = '1' then
			current_state <= inst_fetch;
		elsif clk'event and clk = '1' then 
			case current_state is
				when inst_fetch => 
					current_state <= inst_decode_reg_fetch;
				when inst_decode_reg_fetch => 
					if opcode = "000000" then -- R-type	
						current_state <= execution;
					elsif opcode = "100011" or opcode = "101011" then -- LW/SW
						current_state <= mem_comp;
					elsif opcode = "000100" then -- Beq	
						current_state <= branch_comp;
					elsif opcode = "000010" then -- J-type
						current_state <= jump_comp;
					end if;
				when mem_comp =>	
					if opcode = "100011" then -- LW
						current_state <= mem_r;
					elsif opcode = "101011" then -- SW
						current_state <= mem_w;
					end if;
				when execution => 
					current_state <= r_comp;
				when branch_comp => 
					current_state <= inst_fetch;
				when jump_comp => 
					current_state <= inst_fetch;
				when mem_r => 
					current_state <= write_back;
				when mem_w => 
					current_state <= inst_fetch;
				when r_comp =>
					current_state <= inst_fetch;
				when write_back => 
					current_state <= inst_fetch;
				when others =>
					null;
			end case;
		end if;
	end process;	  
end architecture;